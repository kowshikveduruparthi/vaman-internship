//F =1
module two(x,y,z,a,b,c,d,e,f,g);
  output a,b,c,d,e,f,g;
  input x,y,z;
  //reg F;
   

   not(F,1);  

    /*buf(a,1);
    not(b,1);
    not(c,1);
    buf(d,1);
    buf(e,1);
     buf(f,1);
      buf(g,1);*/
 
endmodule
